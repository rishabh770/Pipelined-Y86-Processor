module sub64_test();

    reg signed [63:0]a;
	reg signed [63:0]b;
    reg signed cin;
    wire signed [63:0]result;
    wire signed overflow;

    sub_64bit dut(.a(a),.b(b),.cin(cin),.result(result),.overflow(overflow));

    initial
    begin
        $dumpfile("sub_out.vcd");
        $dumpvars(0,sub64_test);
        assign a = 64'b0000000000000000000000000000000000000000000000000000000000001111;
        assign b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        assign cin = 1'b0;
        #50;
        assign a = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        assign b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        assign cin = 1'b0;
        #50;
        assign a = 64'b0000100011001001101010010111110010100111101000101001011101011010;
        assign b = 64'b1010101111101010101100101011010110101101101010101010101010101001;
        assign cin = 1'b0;
        #50;
        assign a = 64'b0000000000000000101101001001010110100010000001000100010011101111;
        assign b = 64'b0000000000000000000000000101010100101010010100010101001010101010;
        assign cin = 1'b0;
        #50;
        assign a = 64'b0000001111111010010000000010101111111111000101001111110000000110;
        assign b = 64'b1111111111111111111110010000001001011111100100000001101011110001;
        assign cin = 1'b0;
        #50;
        assign a = 64'b0000000000000000000000000000000000000000100010000000000010001001;
        assign b = 64'b0000000000000000000000000000000000000000000000010010011111111001;
        assign cin = 1'b0;
        #50;
        assign a = 64'b1111111111111111111111111111111111111111111111111110010010000100;
        assign b = 64'b1111111100000001001011111000010010001001010100010000111110010011;
        assign cin = 1'b0;
        #50;
        assign a = 64'b1100010011110101010000000000010010100001111010110110011010111110;
        assign b = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        assign cin = 1'b0;
        #50;

    end
    initial 
    begin
	    $monitor("a=%b\nb=%b\ny=%b\noverflow=%b\n",a,b,result,overflow);
    end

endmodule