module xor_test();

    reg [64:1]a;
	reg [64:1]b;

    wire [64:1]result;

    xor_64bit dut(.a(a),.b(b),.result(result));

    initial
    begin
        $dumpfile("xor_out.vcd");
        $dumpvars(0,xor_test);
        //Case 1
        assign a = 64'b11010011;
        assign b = 64'b11010011;
        #50;
        //Case 2
        assign a = 64'b1111010100100111001010100;
        assign b = 64'b11100110101010011010010011;
        #50;
        //Case 3
        assign a = 64'b0100001001010110010010010111101000100010101001010010101001010011;
        assign b = 64'b1101001010101001100101001001010101010100110100100110010100101010;
        #50;
        //Case 4
        assign a = 64'b1101001001110101001001110011101000100010101001010010101001010011;
        assign b = 64'b1110011011010010001000010001010101010100110100100110010100101010;
        #50;
        //Case 5
        assign a = 64'b1010101110101101011000100010101001010010101001010011;
        assign b = 64'b100010011010101010010101001111011010101010110101010;
        #50;

    end
    initial 
    begin
	    $monitor("a=%b\nb=%b\ny=%b\n",a,b,result);
    end

endmodule