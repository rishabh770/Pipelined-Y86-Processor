module and_test();

    reg [64:1]a;
	reg [64:1]b;

    wire [64:1]result;

    and_64bit dut(.a(a),.b(b),.result(result));

    initial
    begin
        $dumpfile("and_out.vcd");
        $dumpvars(0,and_test);
        assign a = 64'b1001000100010001000100010001000100010001000100010001000100010001;
        assign b = 64'b1110111011101110111011101110111011101110111011101110111011101110;
        #50;
        assign a = 64'b0000000000000000000000000000000000000000000000000000000000001111;
        assign b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        #50;
        assign a = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        assign b = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        #50;
        assign a = 64'b0000100011001001101010010111110010100111101000101001011101011010;
        assign b = 64'b1010101111101010101100101011010110101101101010101010101010101001;
        #50;
        assign a = 64'b0000000000000000101101001001010110100010000001000100010011101111;
        assign b = 64'b0000000000000000000000000101010100101010010100010101001010101010;
        #50;
        assign a = 64'b0000001111111010010000000010101111111111000101001111110000000110;
        assign b = 64'b1111111111111111111110010000001001011111100100000001101011110001;
        #50;
        assign a = 64'b0000000000000000000000000000000000000000100010000000000010001001;
        assign b = 64'b0000000000000000000000000000000000000000000000010010011111111001;
        #50;
        assign a = 64'b1111111111111111111111111111111111111111111111111110010010000100;
        assign b = 64'b1111111100000001001011111000010010001001010100010000111110010011;
        #50;
        assign a = 64'b1100010011110101010000000000010010100001111010110110011010111110;
        assign b = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        #50;
    end
    initial 
    begin
	    $monitor("a=%b\nb=%b\ny=%b\n",a,b,result);
    end

endmodule
